module Sch_Lab407ND(
    );


endmodule
